
class Packet;
    rand bit [2:0] data;
endclass

